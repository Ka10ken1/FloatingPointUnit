// `include "../multree.sv"

module tb_multree;
  reg [57:0] a;
  reg [57:0] b;
  wire [115:0] out;
  multree uut (
    .a(a),
    .b(b),
    .out(out)
  );

  initial begin
    $monitor("Time = %0t | a = %d | b = %d | out = %d", $time, a, b, out);

    a = 58'b00000000000000000000000000000000000000000000000000000001100;
    b = 58'b00000000000000000000000000000000000000000000000000000001100;
    #10;  

    a = 58'b00000000000000000000000000000000000000000000000000000000010;
    b = 58'b00000000000000000000000000000000000000000000000000000000001;
    #10;

    a = 58'b01010101010101010101010101010101010101010101010101010101010;
    b = 58'b01100110011001100110011001100110011001100110011001100110011;
    #10;

  end
endmodule

