// `include "./../lrs.sv"
module tb_lrs;
    reg [6:0] as2;
    reg [54:0] fb2;
    wire [54:0] fb3;

    lrs uut (
        .as2(as2),
        .fb2(fb2),
        .fb3(fb3)
    );

    initial begin
        $display("Time | as2     | fb2                                         | fb3");
        $monitor("%4t | %b      | %b | %b", $time, as2, fb2, fb3);

        as2 = 7'b1010101;
        fb2 = 55'b11011010110111010110111010110111010110111011011010110;  // 55 bits exact
        #10;

        as2 = 7'b0000000;
        fb2 = 55'b10101010101010101010101010101010101010101010101010101;  // 55 bits exact
        #10;

        as2 = 7'b1111111;
        fb2 = 55'b00110011001100110011001100110011001100110011001100110;  // 55 bits exact
        #10;

        as2 = 7'b1011101;
        fb2 = 55'b01010101010101010101010101010101010101010101010101010;  // 55 bits exact
        #10;

        as2 = 7'b0001101;
        fb2 = 55'b11111111111111111111111111111111111111111111111111111;  // 55 bits exact
        #10;
        
        $stop;
    end

endmodule

